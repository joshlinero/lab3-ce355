library IEEE;
use IEEE.std_logic_1164.all;
--Additional standard or custom libraries go here

entity display_divider is
	port(
		--You will replace these with your actual inputs and outputs
		inputs : in std_logic;
		outputs : out std_logic
	 );
end entity display_divider;

architecture structural of display_divider is
--Signals and components go here

begin
--Structural design goes here

end architecture structural;