library IEEE;
use IEEE.std_logic_1164.all; -- Include any additional libraries if needed

package decoder is
    COMPONENT leddcdc
        PORT (
            data_in : in std_logic_vector(3 downto 0);  -- Input port for data
            segments_out : out std_logic_vector(6 downto 0)  -- Output port for segments
        );
    end COMPONENT;
    
    -- Additional components can be declared here if needed in the future

end package decoder;

package body decoder is
    -- Subroutine declarations go here if you have functions or procedures to include
end package body decoder;
